.include p18_cmos_models_tt.inc

.param W = 1u
.param L = 1u
.param Ib = 6.43u

Vdd 0 vdd 1

Ibias_1 vdd ibias_1 4*Ib
Ibias_2 vdd ibias_2 Ib
Ibias_3 vdd ibias_3 Ib
Ibias_4 vdd ibias_4 4*Ib
Iin     vdd iin     7*Ib

*DRAIN GATE SOURCE BASE
mn1     vout        ibias_1     Q1_S    0   NMOS    l = L   w = W
mn2     Q1_S        iin         0       0   NMOS    l = L   w = W
mn3     ibias_1     ibias_2     0       0   NMOS    l = L   w = W
mn4     ibias_2     ibias_2     Q1_S    0   NMOS    l = L   w = W

mn5     iin         ibias_4     Q5_S    0   NMOS    l = L   w = W
mn6     Q5_S        iin         0       0   NMOS    l = L   w = W
mn7     ibias_4     ibias_3     0       0   NMOS    l = L   w = W
mn8     ibias_3     ibias_3     Q5_S    0   NMOS    l = L   w = W

Vout vout 0 0